`include "../00_TESTBED/pseudo_DRAM.sv"
`include "Usertype_OS.sv"

program automatic PATTERN(input clk, INF.PATTERN inf);
import usertype::*;

//================================================================
// parameters & integer
//================================================================
parameter DRAM_p_r = "../00_TESTBED/DRAM/dram.dat";
logic[7:0] golden_DRAM[ ((65536+256*8)-1):(65536+0)];
initial $readmemh(DRAM_p_r, golden_DRAM);
integer gap,lat,y,i;
Error_Msg golden_err;
logic golden_complete;
logic [31:0]golden_info;

//================================================================
// initial
//================================================================
initial begin
	golden_complete = 0;
	golden_info = 0;
	golden_err = No_Err;
	reset_signal_task;
	input_task_output;
	YOU_PASS_task;
	$finish;
end
task input_task_output;begin
	//begin //1
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd162;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd44;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 32'b100110101101100100000100101100;
	golden_err = No_Err;
	tastoutput;
	// 2
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 32'b10011010110110;
	golden_err = No_Err;
	tastoutput;
	// 3
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 15'b110101001111001;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 32'b1001000100101111;
	golden_err = No_Err;
	tastoutput;
	// 4
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd45;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd45;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hca;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	// 5
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd84;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h7670;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//6
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd48;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h67;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//7
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd33;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd25;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	// 8
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he348;
	golden_err = No_Err;
	tastoutput;
	//9
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hde;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd50;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd64;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//10
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd24;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8f;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//11
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h6489;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9124;
	golden_err = No_Err;
	tastoutput;
	//12
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd33;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h7b;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//13
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd45;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd65;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//14
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h68;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd42;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd46;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//15
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h69;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hbb334169;
	golden_err = No_Err;
	tastoutput;
	//16
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd163;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd35;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Out_of_money;
	tastoutput;
	//17
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd24;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd144;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//18
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb8;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h6a9a;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc259;
	golden_err = No_Err;
	tastoutput;
	//19
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd66;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1ae;
	golden_err = No_Err;
	tastoutput;
	//20 //27
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hcc;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h62d9;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf7e1;
	golden_err = No_Err;
	tastoutput;
	//21 //29
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd164;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd12;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd165;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc60c4ca5;
	golden_err = No_Err;
	tastoutput;
	//22 //31
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd18;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd47;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h17a2d22f;
	golden_err = No_Err;
	tastoutput;
	//23 //32
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hda84;
	golden_err = No_Err;
	tastoutput;
	//24 //34
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h7e;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc936967e;
	golden_err = No_Err;
	tastoutput;
	//25 //35
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h6a;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hbfb8486a;
	golden_err = No_Err;
	tastoutput;
	//26 //36
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd27;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h58c7;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h84da;
	golden_err = No_Err;
	tastoutput;
	//27 //37
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd67;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 3;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd38;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h92;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h4ec7e692;
	golden_err = No_Err;
	tastoutput;
	//28 //38
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9fd7;
	golden_err = No_Err;
	tastoutput;
	//29 //39
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'he1b9;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//30 //40
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd87;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd49;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd28;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//31 //41
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h6736;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h8b67;
	golden_err = No_Err;
	tastoutput;
	//32 //43
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hcd;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h864c;
	golden_err = No_Err;
	tastoutput;
	//33 //44
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd48;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd37;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd26;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//34 //45
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h7f;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h2d2e2;
	golden_err = No_Err;
	tastoutput;
	//35 //46
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd86;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h5507;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//36 //47
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd36;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hba;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//37 //48
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb9;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd35;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd68;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//38 //50
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd9;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//39 //53
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h93;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd31;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd49;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc853df31;
	golden_err = No_Err;
	tastoutput;
	//40 //54
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd107;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf6;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//41 //55
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h5abf;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7fa7;
	golden_err = No_Err;
	tastoutput;
	//42 //56
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd27;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h80;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//43 //57
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hbb;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd35;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h91;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//44 //60
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hcf;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd27;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hce;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//45 //61
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd167;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd44;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd168;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//46 //63
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd6;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hde79c6e2;
	golden_err = No_Err;
	tastoutput;
	//47 //64
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9402;
	golden_err = No_Err;
	tastoutput;
	//48 //69
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd11;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd6;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//49 //73
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h6e;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hfd8c;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//50 //74
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd31;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h4da1c41f;
	golden_err = No_Err;
	tastoutput;
	//51 //76
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd169;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3de3e8a9;
	golden_err = No_Err;
	tastoutput;
	//52 //77
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd51;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h6782;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hae72;
	golden_err = No_Err;
	tastoutput;
	//53 //78
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'h2b;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h81;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//54 //84
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd170;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'h1a;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h6f;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//55 //86
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd32;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hefea;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//56 //91
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h5b;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9df3835b;
	golden_err = No_Err;
	tastoutput;
	//57 //92
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h5b;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3c4d7;
	golden_err = No_Err;
	tastoutput;
	//58 //93
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hb490;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//59 //94
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd37;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd52;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//60 //96
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'he5fd;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//61 //97
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h83;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//62 //98
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h96;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd7;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hbe;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h62acc7be;
	golden_err = No_Err;
	tastoutput;
	//63 //99
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h48;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd46;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf8;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//64 //100
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hfa;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h70;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7418;
	golden_err = No_Err;
	tastoutput;
	//65 //101
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he6;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h6aa9c4e6;
	golden_err = No_Err;
	tastoutput;
	//66 //102
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hc2e9;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//67 //103
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he6;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h36cdf;
	golden_err = No_Err;
	tastoutput;
	//68 //108
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd33;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd15;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd34;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7fab4f22;
	golden_err = No_Err;
	tastoutput;
	//69 //110
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hbf;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hb1c5;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he28e;
	golden_err = No_Err;
	tastoutput;
	//70 //112
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h1314;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h8d5e;
	golden_err = No_Err;
	tastoutput;
	//71 //113
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd54;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h8ac4;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//72 //114
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd7;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd14;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//73 //115
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd15;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h6418810f;
	golden_err = No_Err;
	tastoutput;
	//74 //116
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h98;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_ID;
	tastoutput;
	//75 //117
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd92;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5fea855c;
	golden_err = No_Err;
	tastoutput;
	//76 //118
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd35;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb0405323;
	golden_err = No_Err;
	tastoutput;
	//77 //121
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hfb;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd28;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd74;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//78 //123
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h72;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h559e;
	golden_err = No_Err;
	tastoutput;
	//79 //124
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd21;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd55;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//80 //126
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h85;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd53;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h287fd635;
	golden_err = No_Err;
	tastoutput;
	//81 //132
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he9;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h38c2;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hebb9;
	golden_err = No_Err;
	tastoutput;
	//82 //135
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd26;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd75;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he173da4b;
	golden_err = No_Err;
	tastoutput;
	//83 //137
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h73;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hafb5;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//84 //138
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h5f;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd25;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hfd;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//85 //140
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd36;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h70ab;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h8252;
	golden_err = No_Err;
	tastoutput;
	//86 //144
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd6;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h87;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//87 //145
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h517c;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h97df;
	golden_err = No_Err;
	tastoutput;
	//88 //146
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd37;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//89 //147
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h39;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd37;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd17;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//90 //150
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hfe;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h20fd;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf4be;
	golden_err = No_Err;
	tastoutput;
	//91 //151
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd18;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h8b1b;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9bad;
	golden_err = No_Err;
	tastoutput;
	//92 //152
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd38;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//93 //153
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd12;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd77;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//94 //155
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hea;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h900c;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//95 //156
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h6dfd;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he0e1;
	golden_err = No_Err;
	tastoutput;
	//96 //157
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hb01a;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//97 //158
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd46;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd96;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//98 //160
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h5d5;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h2e4b;
	golden_err = No_Err;
	tastoutput;
	//99 //162
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd97;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//100 //163
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h8579;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb3c4;
	golden_err = No_Err;
	tastoutput;
	//101 //164
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd58;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd47;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'heb;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//102 //165
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h85eb83b0;
	golden_err = No_Err;
	tastoutput;
	//103 //166
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h4e;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3b10d;
	golden_err = No_Err;
	tastoutput;
	//104 //167
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h9d;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h30f3e;
	golden_err = No_Err;
	tastoutput;
	//105 //168
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd47;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd174;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//106 //170
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h74;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hca2b;
	golden_err = No_Err;
	tastoutput;
	//107 //171
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd39;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf780;
	golden_err = No_Err;
	tastoutput;
	//108 //172
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h7a47;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'ha20f;
	golden_err = No_Err;
	tastoutput;
	//109 //176
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd44;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd98;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//110 //178
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd27;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd59;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//111 //179
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd9;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//112 //180
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8a;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd6;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//113 //181
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd24;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//114 //182
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd21;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//115 //184
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hed;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd12;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd80;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf83ccc50;
	golden_err = No_Err;
	tastoutput;
	//116 //185
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h9e33;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc304;
	golden_err = No_Err;
	tastoutput;
	//117 //186
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd21;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h9c7;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he5c3;
	golden_err = No_Err;
	tastoutput;
	//118 //187
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd27;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h9e;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//119 //188
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h9f;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd28;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hda;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//120 //190
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h77;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 3;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd45;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd100;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//121 //191
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd33;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8b;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//122 //192
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h4487;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'he489;
	golden_err = No_Err;
	tastoutput;
	//123 //193
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hce275302;
	golden_err = No_Err;
	tastoutput;
	//124 //194
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd48;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h3c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_ID;
	tastoutput;
	//125 //196
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd41;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h78;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3df92;
	golden_err = No_Err;
	tastoutput;
	//126 //197
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd50;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h3d;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//127 //199
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd11;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h39f14bc7;
	golden_err = No_Err;
	tastoutput;
	//128 //200
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd23;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd101;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//129 //201
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd11;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc7;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h2de29;
	golden_err = No_Err;
	tastoutput;
	//130 //204
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hef;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//131 //206
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h79;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd50;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd62;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//132 //207
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd17;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8d;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//133 //209
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd160;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd10;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd82;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//134 //210
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hec;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd24;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hb3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//135 //212
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h2b;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd161;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7ef583a1;
	golden_err = No_Err;
	tastoutput;
	//136 //213
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h66;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd23;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3406c317;
	golden_err = No_Err;
	tastoutput;
	//137 //214
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd34;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc8;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//138 //215
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hde6d;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfd86;
	golden_err = No_Err;
	tastoutput;
	//139 //221
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd26;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//140 //223
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8e;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h3f5d;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'ha065;
	golden_err = No_Err;
	tastoutput;
	//141 //225
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hdb;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd11;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd161;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//142 //226
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd19;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'he5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//143 //230
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h8c9;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hcb8b;
	golden_err = No_Err;
	tastoutput;
	//144 //231
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd48;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd28;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//145 //233
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hcb;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd39;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd54;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Out_of_money;
	tastoutput;
	//146 //235
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd14;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Not_Enough;
	tastoutput;
	//147
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc282c102;
	golden_err = No_Err;
	tastoutput;
	//148
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h397ac101;
	golden_err = No_Err;
	tastoutput;
	//149
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5f40c101;
	golden_err = No_Err;
	tastoutput;
	//150
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc2c8c1c0;
	golden_err = No_Err;
	tastoutput;
	//151
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb30ae803;
	golden_err = No_Err;
	tastoutput;
	//152
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9dc7e801;
	golden_err = No_Err;
	tastoutput;
	//153
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb2ece803;
	golden_err = No_Err;
	tastoutput;
	//154
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9da9e801;
	golden_err = No_Err;
	tastoutput;
	//155
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb2cee803;
	golden_err = No_Err;
	tastoutput;
	//156
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9d8be801;
	golden_err = No_Err;
	tastoutput;
	//157
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb2b0e803;
	golden_err = No_Err;
	tastoutput;
	//158
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9d6de801;
	golden_err = No_Err;
	tastoutput;
	//159
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1e2c103;
	golden_err = No_Err;
	tastoutput;
	//160
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h9d4fc101;
	golden_err = No_Err;
	tastoutput;
	//161
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1748102;
	golden_err = No_Err;
	tastoutput;
	//162
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h395c8101;
	golden_err = No_Err;
	tastoutput;
	//163
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1064102;
	golden_err = No_Err;
	tastoutput;
	//164
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h393e4101;
	golden_err = No_Err;
	tastoutput;
	//165
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e324101;
	golden_err = No_Err;
	tastoutput;
	//166
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc22841c0;
	golden_err = No_Err;
	tastoutput;
	//166
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc228;
	golden_err = No_Err;
	tastoutput;
	//167
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1bac102;
	golden_err = No_Err;
	tastoutput;
	//168
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3920c101;
	golden_err = No_Err;
	tastoutput;
	//169
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb274e88c;
	golden_err = No_Err;
	tastoutput;
	//170
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf019e801;
	golden_err = No_Err;
	tastoutput;
	//171
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb26ae88c;
	golden_err = No_Err;
	tastoutput;
	//172
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hefd3e801;
	golden_err = No_Err;
	tastoutput;
	//173
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb260e88c;
	golden_err = No_Err;
	tastoutput;
	//174
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hefa1e801;
	golden_err = No_Err;
	tastoutput;
	//175
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb256e88c;
	golden_err = No_Err;
	tastoutput;
	//176
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hef6fe801;
	golden_err = No_Err;
	tastoutput;
	//177
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb24ce88c;
	golden_err = No_Err;
	tastoutput;
	//178
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hef3de801;
	golden_err = No_Err;
	tastoutput;
	//179
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb242e88c;
	golden_err = No_Err;
	tastoutput;
	//180
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hef0be801;
	golden_err = No_Err;
	tastoutput;
	//181
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hd77d5401;
	golden_err = No_Err;
	tastoutput;
	//182
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1d8548c;
	golden_err = No_Err;
	tastoutput;
	//183
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hd75f5401;
	golden_err = No_Err;
	tastoutput;
	//184
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hc1ce548c;
	golden_err = No_Err;
	tastoutput;
	//185
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hb224e88c;
	golden_err = No_Err;
	tastoutput;
	//186
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h8c;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'heeb1e801;
	golden_err = No_Err;
	tastoutput;
	//187
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa4a9ec0;
	golden_err = No_Err;
	tastoutput;
	//188
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5f189e01;
	golden_err = No_Err;
	tastoutput;
	//189
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa409ec0;
	golden_err = No_Err;
	tastoutput;
	//190
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5ee69e01;
	golden_err = No_Err;
	tastoutput;
	//191
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa369ec0;
	golden_err = No_Err;
	tastoutput;
	//192
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5eb49e01;
	golden_err = No_Err;
	tastoutput;
	//193
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa2c9ec0;
	golden_err = No_Err;
	tastoutput;
	//194
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e829e01;
	golden_err = No_Err;
	tastoutput;
	//195
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa229ec0;
	golden_err = No_Err;
	tastoutput;
	//196
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e649e01;
	golden_err = No_Err;
	tastoutput;
	//197
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa189ec0;
	golden_err = No_Err;
	tastoutput;
	//198
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e469e01;
	golden_err = No_Err;
	tastoutput;
	//199
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa0e9ec0;
	golden_err = No_Err;
	tastoutput;
	//200
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e289e01;
	golden_err = No_Err;
	tastoutput;
	//201
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'haa049ec0;
	golden_err = No_Err;
	tastoutput;
	//202
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e0a9e01;
	golden_err = No_Err;
	tastoutput;
	//203
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'ha9fa9ec0;
	golden_err = No_Err;
	tastoutput;
	//204
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd30;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'h1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5e009e01;
	golden_err = No_Err;
	tastoutput;
	//205
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h494e6802;
	golden_err = No_Err;
	tastoutput;
	//206
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//206
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h491c6802;
	golden_err = No_Err;
	tastoutput;
	//207
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//208
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h48ea6802;
	golden_err = No_Err;
	tastoutput;
	//209
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//210
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h48cc6802;
	golden_err = No_Err;
	tastoutput;
	//211
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//212
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h48ae6802;
	golden_err = No_Err;
	tastoutput;
	//213
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//214
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd16;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h48a46802;
	golden_err = No_Err;
	tastoutput;
	//215
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd40;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h7259;
	golden_err = No_Err;
	tastoutput;
	//216
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'h3e90;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfffa;
	golden_err = No_Err;
	tastoutput;
	//217
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h389ec101;
	golden_err = No_Err;
	tastoutput;
	//218
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hffff;
	golden_err = No_Err;
	tastoutput;
	//219
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hff91c102;
	golden_err = No_Err;
	tastoutput;
	//220
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h381c8101;
	golden_err = No_Err;
	tastoutput;
	//221
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hffff;
	golden_err = No_Err;
	tastoutput;
	//222
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hff2d8102;
	golden_err = No_Err;
	tastoutput;
	//224
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h379a4101;
	golden_err = No_Err;
	tastoutput;
	//225
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hffff;
	golden_err = No_Err;
	tastoutput;
	//226
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfec94102;
	golden_err = No_Err;
	tastoutput;
	//227
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'ha3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd35;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Out_of_money;
	tastoutput;
	//228
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hd556f3;
	golden_err = No_Err;
	tastoutput;
	//229
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Out_of_money;
	tastoutput;
	//230
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Out_of_money;
	tastoutput;
	//231
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd22;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h239f;
	golden_err = No_Err;
	tastoutput;
	//232
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h27df45f3;
	golden_err = No_Err;
	tastoutput;
	//233
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//234
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h27ad45f3;
	golden_err = No_Err;
	tastoutput;
	//235
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//236
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h277b45f3;
	golden_err = No_Err;
	tastoutput;
	//237
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//238
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h23c548f3;
	golden_err = No_Err;
	tastoutput;
	//239
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//240
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h158354f3;
	golden_err = No_Err;
	tastoutput;
	//241
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//242
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h155154f3;
	golden_err = No_Err;
	tastoutput;
	//243
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd20;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//242
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd9;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h221749f3;
	golden_err = No_Err;
	tastoutput;
	//243
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd9;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hf3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f0b0;
	golden_err = No_Err;
	tastoutput;
	//244
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfd934102;
	golden_err = No_Err;
	tastoutput;
	//245
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_ID;
	tastoutput;
	//246
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hebad4105;
	golden_err = No_Err;
	tastoutput;
	//247
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_Num;
	tastoutput;
	//248
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_Item;
	tastoutput;
	//249
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3beff;
	golden_err = No_Err;
	tastoutput;
	//250
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfc5d4102;
	golden_err = No_Err;
	tastoutput;
	//251
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//252
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd60;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//253
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'heb8f4102;
	golden_err = No_Err;
	tastoutput;
	//254
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	//255
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfb274102;
	golden_err = No_Err;
	tastoutput;
	//256
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hffff;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//257
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd3;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_ID;
	tastoutput;
	//258
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_Num;
	tastoutput;
	//259
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_Item;
	tastoutput;
	//260
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1f604;
	golden_err = No_Err;
	tastoutput;
	//261
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hea454105;
	golden_err = No_Err;
	tastoutput;
	//262
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'hffff;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wallet_is_Full;
	tastoutput;
	//263
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd10;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd15;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1802410f;
	golden_err = No_Err;
	tastoutput;
	//264
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h1802;
	golden_err = No_Err;
	tastoutput;
	//265
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd60;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd10;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = INV_Full;
	tastoutput;
	//266
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd5;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3ceff;
	golden_err = No_Err;
	tastoutput;
	//267
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hfb1d4102;
	golden_err = No_Err;
	tastoutput;
	//268
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h3c2c4101;
	golden_err = No_Err;
	tastoutput;
	//269
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd8;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 0;
	golden_info = 0;
	golden_err = Wrong_act;
	tastoutput;
	for(i=0;i<256;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = i;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'hffff;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
	end
	for(i=0;i<256;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = i;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'hffff;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
	end
	for(i=0;i<20;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'd45;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.item_valid = 1;
		inf.D = 'd2;
		@(negedge clk);
		inf.item_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.num_valid = 1;
		inf.D = 'd16;
		@(negedge clk);
		inf.num_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'd65;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = INV_Not_Enough;
		tastoutput;
		///
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'd163;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.item_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.item_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.num_valid = 1;
		inf.D = 'd35;
		@(negedge clk);
		inf.num_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'hf3;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Out_of_money;
		tastoutput;
	end
	//////
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'hc0;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.item_valid = 1;
	inf.D = 'd2;
	@(negedge clk);
	inf.item_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.num_valid = 1;
	inf.D = 'd1;
	@(negedge clk);
	inf.num_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.id_valid = 1;
	inf.D = 'd15;
	@(negedge clk);
	inf.id_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'h5d2e810f;
	golden_err = No_Err;
	tastoutput;
	///////
	for(i=0;i<20;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd8;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.item_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.item_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.num_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.num_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'h98;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wrong_ID;
		tastoutput;
	end	
	for(i=0;i<20;i=i+1)begin
		////73 //115
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd8;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.item_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.item_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.num_valid = 1;
		inf.D = 'd3;
		@(negedge clk);
		inf.num_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'd15;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wrong_Num;
		tastoutput;
	end
	for(i=0;i<20;i=i+1)begin
		////73 //115
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd8;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.item_valid = 1;
		inf.D = 'd3;
		@(negedge clk);
		inf.item_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.num_valid = 1;
		inf.D = 'd1;
		@(negedge clk);
		inf.num_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.id_valid = 1;
		inf.D = 'd15;
		@(negedge clk);
		inf.id_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wrong_Item;
		tastoutput;
	end
	//////
	gap = $urandom_range(3,8);
	repeat(gap)@(negedge clk);
	inf.act_valid = 1;
	inf.D = 'd4;
	@(negedge clk);
	inf.act_valid = 0;
	inf.D = 'dx;
	gap = $urandom_range(1,4);
	repeat(gap)@(negedge clk);
	inf.amnt_valid = 1;
	inf.D = 'd40000;
	@(negedge clk);
	inf.amnt_valid = 0;
	inf.D = 'dx;
	golden_complete = 1;
	golden_info = 'hf96e;
	golden_err = No_Err;
	tastoutput;
	for(i=0;i<20;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'd10000;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
		///
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'd20000;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
		////gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'd40000;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
		///
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd4;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		gap = $urandom_range(1,4);
		repeat(gap)@(negedge clk);
		inf.amnt_valid = 1;
		inf.D = 'd50000;
		@(negedge clk);
		inf.amnt_valid = 0;
		inf.D = 'dx;
		golden_complete = 0;
		golden_info = 0;
		golden_err = Wallet_is_Full;
		tastoutput;
	end
	for(i=0;i<100;i=i+1)begin
		gap = $urandom_range(3,8);
		repeat(gap)@(negedge clk);
		inf.act_valid = 1;
		inf.D = 'd2;
		@(negedge clk);
		inf.act_valid = 0;
		inf.D = 'dx;
		golden_complete = 1;
		golden_info = 'hf96e;
		golden_err = No_Err;
		tastoutput;
	end
end endtask
task tastoutput;begin
	wait_OUT_VALID;
	y=0;
	while(inf.out_valid===1)begin
		if(inf.complete !== golden_complete || inf.out_info!== golden_info|| inf.err_msg!==golden_err)begin
			$display ("Wrong Answer");
			$finish;
		end
		@(negedge clk);	
		y=y+1;
	end	 	
end endtask
task wait_OUT_VALID; begin
  lat = -1;
  while(inf.out_valid!==1) begin
	lat = lat + 1;
	if(lat == 10000) begin
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");
		$display ("                                                                        FAIL!                                                               ");
		$display ("                                                     The execution latency are over 10000   cycles                                            ");
		$display ("--------------------------------------------------------------------------------------------------------------------------------------------");

		repeat(2)@(negedge clk);
		$finish;
	end
	@(negedge clk);
  end
end endtask
task reset_signal_task; begin 
	inf.rst_n = 1;
    #(0.5);   inf.rst_n = 0;
	#(2.0);
	inf.id_valid = 0;
	inf.act_valid = 0;
	inf.num_valid = 0;
	inf.item_valid = 0;
	inf.amnt_valid = 0;
	inf.D = 'dx;
	#(10);   inf.rst_n=1;
end endtask
task YOU_PASS_task;begin

$display ("----------------------------------------------------------------------------------------------------------------------");
$display ("                                                  Congratulations!                						            ");
$display ("                                           You have passed all patterns!          						            ");
$display ("----------------------------------------------------------------------------------------------------------------------");
end endtask
endprogram
